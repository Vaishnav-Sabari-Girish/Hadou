//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025-10-10 04:39:29 UTC
// Design Name: NOT_GATE
// Module Name: NOT_GATE
// Project Name: NOT_GATE
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module NOT_GATE (
  input a,b,
  output c
);

and a1(c, a, b);

endmodule
