`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025-10-09 17:32:23 UTC
// Design Name: Test_Verilog
// Module Name: Test_Verilog
// Project Name: Test_Verilog
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module Test_Verilog (
  input a, b,
  output c
);

assign c = a & b;

endmodule
